* C:\Users\DELL\eSim-Workspace\akhil_full_adder\akhil_full_adder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/4/2022 9:34:09 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ akhil_full_adder		
U5  A B Cin Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ adc_bridge_3		
U6  Net-_U1-Pad4_ Net-_U1-Pad5_ Sum Carry dac_bridge_2		
v3  Cin GND pulse		
v2  B GND pulse		
v1  A GND pulse		
U7  Sum plot_v1		
U8  Carry plot_v1		
U2  A plot_v1		
U3  B plot_v1		
U4  Cin plot_v1		

.end
